* RC Filter
V1 inp 0 dc 0 ac 1
R1 inp out 1k
C1 out 0 1n

.ac dec 10 1 1G
.print ac all
.end
