.title rcfiltertb_r_1k_c_1_0000000000000000622815914577798564188970686927859787829220294952392578125n
.option savecurrents
vi0 vss 0 dc 0
vi1 inp vss dc 0.0e0 ac 1.0e0 0.0e0
ri2 inp out r=1.0e3
ci3 out vss c=1.0000000000000000622815914577798564188970686927859787829220294952392578125e-9
.end
